use library IEEE.std_logic_1164.all;

entity reading_tools is
    port (
        
    )